module booth (
    input  wire        clk  ,
	input  wire        rst_n,
	input  wire [15:0] x    ,
	input  wire [15:0] y    ,
	input  wire        start,
	output  reg  [31:0] z    ,
	output wire        busy 
);

// A����+x
reg  [31:0] A;
// B����-x
reg    [31:0] B;
reg[4:0] cnt;
// CΪ���������չ
integer C=32'h8000_0000;



reg mb=0;

assign busy=mb;

// ��������״̬����busy����ģ��
always @(posedge clk or negedge rst_n) begin
	
	if(!rst_n)
// �����ת״̬����ʼ��
	begin
		cnt<=5'h0;
		mb<=0;

	end
else if(start==1'b1)
// ����start�������г�ʼ̬�����⴦��
	begin
		mb <=1'b1;
		cnt<=5'd1;
	end
	
// ������������ cnt!=0
else

begin	
// cnt 17��ʱ�򵽴����״̬��ֹͣ����
	if(cnt==5'd17)
	begin
	cnt<=0;
	mb<=0;
	end
// ����״̬������ÿ������+1
	else if (cnt!=0)
	begin
	cnt<=cnt+1;
	end
end
end


// �������ݿ���ģ��
always@(posedge clk or negedge rst_n)
begin
// ��λ����
if(!rst_n)
	begin
		A<=0;
		B<=0;
		z<=0;

	end
	
// ����start
else  if(start==1'b1)
	// �������ݣ�ֱ�����뵽���ԼӼ��ĸ�λ���������ֱ�Ӽ���ʹ��
	begin
		A[31:16] <= x;
		A[15:0]<=16'b0;
		B[31:16] <= -x;
		B[15:0]<=16'b0;
		z[15:0]<=y;
		z[31:16]<=16'b0;
	end
// ��������״̬
else 
    begin
	case(cnt)
	// ��״̬
		5'd0:begin
		end
	// ��һ�������жϼӼ�
		5'd1:begin
		case(z[0])
			1'b1: z[31:0] <= z+B[31:0];
			1'b0: z[31:0] <= z;
		endcase
		end
	// ����״̬���⴦��
		5'd17:begin
		  z[31:0] <=(z[31]==1)?((z>>1)+C):  (z>>1);
		end
	// ����Ĭ�ϼ���״̬
		default:
			begin
			case(z[1:0])
			2'b00:
			begin
				z[31:0] <=(z[31]==1)?((z>>1)+C): (z>>1);
			end
			2'b01: 
			begin
				z[31:0] <= (z[31]==1)?((z>>1)+C+A): (z>>1)+A;
			end
			2'b10: 
			begin
				z[31:0] <=(z[31]==1)?((z>>1)+C+B):  (z>>1)+B;
			end
			2'b11:
			begin
				z[31:0] <=(z[31]==1)?((z>>1)+C):  (z>>1);
			end
		endcase
			end
		
	endcase
	end

end

endmodule